* ADG408 SPICE Macro-model    
* Description: Converter                                        
* Generic Desc: 15 V, 8 Channel  Analog mux
* Developed by: JOM / ADSC
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (10/1995) - This model was setup with typical leakage currents at +25C for ADG408 
* Copyright 1995, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*
* Parameters modeled include:
*
* END Notes
*
* Node assignments
* 4 - S1, 5 - S2, 6 - S3, 7 - S4, 12 - S5, 11 - S6, 10 - S7
* 9 - S8, 15 - A2, 16 - A1, 1 - A0, 2 - EN
* 8 - D, 13 - VDD, 14 - GND, 3 - VSS
*                    
.SUBCKT ADG408 4 5 6 7 12 11 10 9 15 16 1 2 8 13 14 3
*
* DEMUX SWITCHES (S1-8 ---> D)
*
*     First Section is for control line A0
*
E_A0_2	  200 14   1 14    1
E_A0_1     30 40 201 40   -1
R_A0_1    200 201         1000
C_A0_X2   201 14          100E-12

V_AX_1     40  14          1.6

S_A0_8      9 34 201 14   Sdemux
S_A0_7     10 34 30  14   Sdemux		
S_A0_6     11 33 201 14   Sdemux
S_A0_5     12 33 30  14   Sdemux
S_A0_4      7 32 201 14   Sdemux
S_A0_3      6 32 30  14   Sdemux
S_A0_2      5 31 201 14   Sdemux
S_A0_1      4 31 30  14   Sdemux

C_A0_X1     1 14          4E-12
C_A0_D      1 39          4E-12

*          Input capacitances

C_A0_1      4  14         8E-12
C_A0_2      5  14         8E-12
C_A0_3      6  14	  8E-12
C_A0_4      7  14         8E-12
C_A0_5     12  14         8E-12
C_A0_6     11  14         8E-12
C_A0_7     10  14         8E-12
C_A0_8      9  14         8E-12

C_D_1       8  14         80E-12

*
*	Leakage Current (SX and D ON only) 
*

R_ON_S1     4 500    1.5E12
R_ON_S2	    5 500    1.5E12
R_ON_S3     6 500    1.5E12
R_ON_S4     7 500    1.5E12
R_ON_S5    12 500    1.5E12
R_ON_S6    11 500    1.5E12
R_ON_S7    10 500    1.5E12
R_ON_S8     9 500    1.5E12

SLEAK_ON_D  8 500    8 500  SLEAK
ILEAK_ON_D  8 500    10E-12 		  
*
*	Leakage Current (SX OFF only)
*
*	Leakage Current (D OFF only)
*

S_OFF_D     8  58 80 14	  Sdemux
R_OFF_D    58  14         1E12 
G_OFF_D     8  14 58 14   0.75E-12

*C_OFF_D     58  14                0E-12   
*
*     Second Section is for control line A1
*

E_A1_2	  170 14 16  14    1
E_A1_1     41 40 171 40   -1
R_A1_1    170 171         1000
C_A1_X2   171 14          100E-12

S_A1_4     34 42 171 14     Sdemux
S_A1_3     33 42 41  14     Sdemux
S_A1_2     32 43 171 14    Sdemux
S_A1_1     31 43 41  14    Sdemux

C_A1_X     16 14           4E-12
C_A1_D     16 39           4E-12

*
*     Third Section is for control line A2
*

E_A2_2	  160  14  15  14  1
E_A2_1     46  40 161  40  -1
R_A2_1    160 161          1000
C_A2_X2   161  14          100E-12

S_A2_2     42 39 161 14    Sdemux
S_A2_1     43 39  46 14    Sdemux

C_A2_X     15 14           4E-12
C_A2_D     15 39           4E-12

*
*     Main Series Switch combination
*
*

V_1_A     419   14  15
V_1_B     420   14  -15
V_1_C     421   13  -1        ;sets pos main offset
V_1_D     422    3  2		;sets neg main offset



R_1_C      39   0         1E13
S_1_A     425  39 420  73 SNCM
R_1_A     412 425         29		;sets neg at max d
S_1_B     426  39 419  73 SPCM
R_1_B      73 426         50            ;sets pos at max d
S_1_C      73 412 611  14 SMAINP
S_1_D     412 411  14 612 SMAINN
E_1_E     611  14         VALUE = {(10*V(73,500))/(V(421,500)+0.005)}
E_1_F     612  14         VALUE = {(10*V(73,500))/(V(500,422)+0.005)}
S_1_G     411  39  99   3 SBASE

*
*	Voltage Clamp 
*

D_1_POS     39  13          DClamp  .001
G_1_POS     39  13  39  13  -1E-12
D_2_NEG      3  39          DClamp  .001
G_2_NEG      3  39   3  39  1E-12

*
*     Enable Switch section
*

S_EN_1     73  8  2  14    Sdemux
C_EN_1      2  8           4.2E-12  ; SETS CHARGE INJECTION 

*     Invert Enable Switch section

E_EN0_1     80  14 2 82    -2
V_EN0_1	    82  14          2.5

*
*     Power Supply Current Correction
*

I_PS_1     13  14           80E-6
I_PS_2     14   3           0.0001E-6
E_PS_1     99  14  13  14   1
E_PS_2    500   3  13   3   .5

*
*	Crosstalk 
*

RXT_1      4 52           1E13
RXT_2      5 52           1E13
RXT_3      6 52           1E13
RXT_4      7 52           1E13
RXT_5     12 52           1E13
RXT_6     11 52           1E13
RXT_7     10 52           1E13
RXT_8      9 52           1E13

CXT_1      4 52           1E-12
CXT_2      5 52           1E-12
CXT_3      6 52           1E-12
CXT_4      7 52           1E-12
CXT_5     12 52           1E-12
CXT_6     11 52           1E-12
CXT_7     10 52           1E-12
CXT_8      9 52           1E-12
*
*	OFF Isolation
*
COI_1      4  8           1E-13
COI_2      5  8           1E-13
COI_3      6  8           1E-13
COI_4      7  8           1E-13
COI_5     12  8           1E-13
COI_6     11  8           1E-13
COI_7     10  8           1E-13
COI_8      9  8           1E-13

ROI_1        4 1901         1.6E9
COI_1A    1901    8         10E-12
ROI_2        5 1902         1.6E9
COI_2A    1902    8         10E-12
ROI_3        6 1903         1.6E9
COI_3A    1903    8         10E-12
ROI_4        7 1904         1.6E9
COI_4A    1904    8         10E-12
ROI_5       12 1905         1.6E9
COI_5A    1905    8         10E-12
ROI_6       11 1906         1.6E9
COI_6A    1906    8         10E-12
ROI_7       10 1907         1.6E9
COI_7A    1907    8         10E-12
ROI_8        9 1908         1.6E9
COI_8A    1908    8         10E-12
*
* MODELS USED
*
.MODEL SNCM  VSWITCH (RON=1 ROFF=400001 VON=18 VOFF=-60)
.MODEL SPCM  VSWITCH (RON=450000 ROFF=1 VON=50 VOFF=-13.5)
.MODEL SBASE VSWITCH (RON=27 ROFF=1400 VON=28 VOFF=-10)
.MODEL SMAINP VSWITCH (RON=250001 ROFF=12 VON=24.5 VOFF=0)
.MODEL SMAINN VSWITCH (RON=250001 ROFF=6 VON=24.5 VOFF=0)
.MODEL Sdemux VSWITCH (RON=1 ROFF=1E12 VON=2.0 VOFF=1.4)
.MODEL DClamp D(IS=1E-15 IBV=1E-13 CJO=1E-12)
.MODEL SLEAK VSWITCH (RON=750E9 ROFF=150E9 VON=-15 VOFF=15)
.PARAM GMIN=1E-14
.ENDS ADG408


